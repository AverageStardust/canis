module top (
    output USBPU,
    output PIN_10,
    output PIN_11
);
    assign USBPU = 0;
    assign PIN_10 = 1;
    assign PIN_11 = 0;
endmodule
